CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
420 340 30 100 10
189 83 1534 801
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
3 4 0.208914 0.148699
357 179 470 276
42991634 0
0
6 Title:
5 Name:
0
0
0
52
13 Logic Switch~
5 611 1041 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4116 0 0
2
5.89916e-315 0
0
13 Logic Switch~
5 156 347 0 1 11
0 30
0
0 0 21360 270
2 0V
-6 -21 8 -13
6 chaveC
-20 -31 22 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8776 0 0
2
5.89916e-315 5.26354e-315
0
13 Logic Switch~
5 93 349 0 10 11
0 50 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
6 chaveB
-20 -31 22 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4460 0 0
2
5.89916e-315 5.30499e-315
0
13 Logic Switch~
5 39 347 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
6 chaveA
-20 -31 22 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7489 0 0
2
5.89916e-315 5.32571e-315
0
13 Logic Switch~
5 543 464 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3231 0 0
2
5.89916e-315 5.34643e-315
0
13 Logic Switch~
5 505 464 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-2 -31 5 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7402 0 0
2
5.89916e-315 5.3568e-315
0
9 2-In AND~
219 1290 879 0 3 22
0 3 4 2
0
0 0 624 90
6 74LS08
-21 -24 21 -16
4 U18B
17 -5 45 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
5368 0 0
2
43790.9 0
0
9 2-In AND~
219 1084 1021 0 3 22
0 6 4 7
0
0 0 624 90
6 74LS08
-21 -24 21 -16
4 U18A
17 -5 45 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
7521 0 0
2
43790.9 1
0
8 3-In OR~
219 946 1746 0 4 22
0 14 13 12 3
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 15 0
1 U
8969 0 0
2
43790.9 2
0
9 2-In AND~
219 812 1819 0 3 22
0 11 15 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
8446 0 0
2
43790.9 3
0
9 2-In AND~
219 810 1746 0 3 22
0 10 15 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
4395 0 0
2
43790.9 4
0
9 2-In AND~
219 810 1678 0 3 22
0 10 11 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U16B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
3940 0 0
2
43790.9 5
0
9 2-In XOR~
219 921 1520 0 3 22
0 9 8 6
0
0 0 624 0
6 74LS86
-21 -24 21 -16
4 U17A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
7738 0 0
2
43790.9 6
0
9 2-In XOR~
219 799 1580 0 3 22
0 11 10 8
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
8575 0 0
2
43790.9 7
0
9 Inverter~
13 724 1538 0 2 22
0 9 15
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
5935 0 0
2
43790.9 8
0
8 2-In OR~
219 1253 790 0 3 22
0 16 2 5
0
0 0 624 90
6 74LS32
-21 -24 21 -16
3 U2C
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
7874 0 0
2
43790.9 9
0
9 2-In AND~
219 1234 923 0 3 22
0 18 17 16
0
0 0 624 90
6 74LS08
-21 -24 21 -16
4 U16A
17 -5 45 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
3791 0 0
2
43790.9 10
0
9 2-In AND~
219 961 907 0 3 22
0 20 18 19
0
0 0 624 90
6 74LS08
-21 -24 21 -16
3 U1D
16 -5 37 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
6882 0 0
2
43790.9 11
0
8 3-In OR~
219 876 1254 0 4 22
0 23 22 21 17
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 15 0
1 U
9189 0 0
2
43790.9 12
0
9 2-In AND~
219 753 1351 0 3 22
0 11 9 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
4194 0 0
2
43790.9 13
0
9 2-In AND~
219 752 1272 0 3 22
0 10 9 22
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-32 -27 -11 -19
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
6368 0 0
2
43790.9 14
0
9 2-In AND~
219 749 1202 0 3 22
0 11 10 23
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
7744 0 0
2
43790.9 15
0
9 2-In XOR~
219 856 1068 0 3 22
0 9 24 20
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
9543 0 0
2
43790.9 16
0
9 2-In XOR~
219 737 1089 0 3 22
0 11 10 24
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U5B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
322 0 0
2
43790.9 17
0
8 2-In OR~
219 1074 675 0 3 22
0 26 25 51
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
3329 0 0
2
5.89916e-315 5.36716e-315
0
8 4-In OR~
219 983 746 0 5 22
0 46 48 19 7 25
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U4B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
8980 0 0
2
5.89916e-315 5.37752e-315
0
8 4-In OR~
219 993 550 0 5 22
0 35 38 41 43 26
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
461 0 0
2
5.89916e-315 5.38788e-315
0
9 2-In NOR~
219 624 777 0 3 22
0 9 10 28
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 NOR
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
9339 0 0
2
5.89916e-315 5.39306e-315
0
10 2-In XNOR~
219 615 927 0 3 22
0 10 9 29
0
0 0 624 0
4 4077
-7 -24 21 -16
4 XNOR
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 13 0
1 U
5483 0 0
2
5.89916e-315 5.39824e-315
0
14 Logic Display~
6 1256 730 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 COUT
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8913 0 0
2
5.89916e-315 5.40342e-315
0
14 Logic Display~
6 1315 631 0 1 2
10 51
0
0 0 53856 0
6 100MEG
3 -16 45 -8
5 SAIDA
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
363 0 0
2
5.89916e-315 5.4086e-315
0
5 7415~
219 283 1247 0 4 22
0 30 50 49 4
0
0 0 624 0
6 74LS15
-21 -28 21 -20
7 ConSUBT
-39 -27 10 -19
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 9 0
1 U
3896 0 0
2
5.89916e-315 5.41378e-315
0
5 7415~
219 282 1122 0 4 22
0 31 50 49 18
0
0 0 624 0
6 74LS15
-21 -28 21 -20
7 ConSOMA
-26 -25 23 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 9 0
1 U
5231 0 0
2
5.89916e-315 5.41896e-315
0
5 7415~
219 286 909 0 4 22
0 30 32 49 47
0
0 0 624 0
6 74LS15
-21 -28 21 -20
7 ConXNOR
-26 -25 23 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 8 0
1 U
6725 0 0
2
5.89916e-315 5.42414e-315
0
5 7415~
219 296 832 0 4 22
0 31 32 49 45
0
0 0 624 0
6 74LS15
-21 -28 21 -20
6 ConXOR
-22 -25 20 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 8 0
1 U
5409 0 0
2
5.89916e-315 5.42933e-315
0
5 7415~
219 295 742 0 4 22
0 30 50 27 42
0
0 0 624 0
6 74LS15
-21 -28 21 -20
6 ConNOR
-22 -25 20 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 8 0
1 U
9227 0 0
2
5.89916e-315 5.43192e-315
0
5 7415~
219 295 664 0 4 22
0 31 50 27 40
0
0 0 624 0
6 74LS15
-21 -28 21 -20
5 ConOR
-18 -25 17 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 7 0
1 U
895 0 0
2
5.89916e-315 5.43451e-315
0
5 7415~
219 297 574 0 4 22
0 30 32 27 37
0
0 0 624 0
6 74LS15
-21 -28 21 -20
7 ConNAND
-26 -26 23 -18
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 7 0
1 U
6121 0 0
2
5.89916e-315 5.4371e-315
0
5 7415~
219 292 506 0 4 22
0 31 32 27 34
0
0 0 624 0
6 74LS15
-21 -28 21 -20
6 ConAND
-26 -30 16 -22
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 7 0
1 U
3291 0 0
2
5.89916e-315 5.43969e-315
0
9 Inverter~
13 218 404 0 2 22
0 30 31
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
8348 0 0
2
5.89916e-315 5.44228e-315
0
9 Inverter~
13 129 401 0 2 22
0 50 32
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
3351 0 0
2
5.89916e-315 5.44487e-315
0
9 Inverter~
13 64 399 0 2 22
0 49 27
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
988 0 0
2
5.89916e-315 5.44746e-315
0
9 2-In AND~
219 733 935 0 3 22
0 29 47 48
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3507 0 0
2
5.89916e-315 5.45005e-315
0
9 2-In AND~
219 737 861 0 3 22
0 44 45 46
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
5175 0 0
2
5.89916e-315 5.45264e-315
0
9 2-In XOR~
219 615 852 0 3 22
0 10 9 44
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 XOR
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3568 0 0
2
5.89916e-315 5.45523e-315
0
9 2-In AND~
219 740 787 0 3 22
0 28 42 43
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
4348 0 0
2
5.89916e-315 5.45782e-315
0
9 2-In AND~
219 747 708 0 3 22
0 39 40 41
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3453 0 0
2
5.89916e-315 5.46041e-315
0
10 2-In NAND~
219 632 599 0 3 22
0 9 10 36
0
0 0 624 0
6 74LS00
-14 -24 28 -16
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
534 0 0
2
5.89916e-315 5.463e-315
0
8 2-In OR~
219 624 699 0 3 22
0 9 10 39
0
0 0 624 0
6 74LS32
-21 -24 21 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7640 0 0
2
5.89916e-315 5.46559e-315
0
9 2-In AND~
219 734 607 0 3 22
0 36 37 38
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U13D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4129 0 0
2
5.89916e-315 5.46818e-315
0
9 2-In AND~
219 724 509 0 3 22
0 33 34 35
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U13B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
6804 0 0
2
5.89916e-315 5.47077e-315
0
9 2-In AND~
219 635 499 0 3 22
0 9 10 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 AND
-13 -29 8 -21
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3264 0 0
2
5.89916e-315 5.47207e-315
0
111
2 3 2 0 0 4224 0 16 7 0 0 3
1265 806
1265 855
1289 855
4 1 3 0 0 8320 0 9 7 0 0 3
979 1746
1280 1746
1280 900
0 2 4 0 0 8320 0 0 7 5 0 4
342 1222
342 1299
1298 1299
1298 900
3 1 5 0 0 4224 0 16 30 0 0 4
1256 760
1256 745
1256 745
1256 748
4 2 4 0 0 0 0 32 8 0 0 4
304 1247
304 1222
1092 1222
1092 1042
3 1 6 0 0 8320 0 13 8 0 0 3
954 1520
1074 1520
1074 1042
4 3 7 0 0 12416 0 26 8 0 0 4
966 760
966 850
1083 850
1083 997
2 3 8 0 0 8320 0 13 14 0 0 4
905 1529
881 1529
881 1580
832 1580
0 1 9 0 0 4096 0 0 13 111 0 4
505 1493
880 1493
880 1511
905 1511
2 0 10 0 0 4096 0 14 0 0 110 2
783 1589
543 1589
1 0 11 0 0 4096 0 14 0 0 100 2
783 1571
610 1571
3 3 12 0 0 4224 0 10 9 0 0 3
833 1819
933 1819
933 1755
2 3 13 0 0 4224 0 9 11 0 0 2
934 1746
831 1746
3 1 14 0 0 4224 0 12 9 0 0 3
831 1678
933 1678
933 1737
1 0 10 0 0 4096 0 12 0 0 110 2
786 1669
543 1669
0 1 10 0 0 0 0 0 11 110 0 3
543 1721
786 1721
786 1737
2 0 15 0 0 4096 0 11 0 0 20 2
786 1755
727 1755
2 0 11 0 0 4096 0 12 0 0 100 2
786 1687
610 1687
1 0 11 0 0 4096 0 10 0 0 100 2
788 1810
610 1810
2 2 15 0 0 4224 0 15 10 0 0 3
727 1556
727 1828
788 1828
0 1 9 0 0 0 0 0 15 111 0 3
505 1508
727 1508
727 1520
3 1 16 0 0 8320 0 17 16 0 0 4
1233 899
1244 899
1244 806
1247 806
4 2 17 0 0 4224 0 19 17 0 0 3
909 1254
1242 1254
1242 944
0 1 18 0 0 8320 0 0 17 27 0 4
354 1122
354 1170
1224 1170
1224 944
3 3 19 0 0 8320 0 26 18 0 0 4
966 751
911 751
911 883
960 883
3 1 20 0 0 8320 0 23 18 0 0 3
889 1068
951 1068
951 928
4 2 18 0 0 0 0 33 18 0 0 4
303 1122
974 1122
974 928
969 928
3 3 21 0 0 8320 0 20 19 0 0 4
774 1351
859 1351
859 1263
863 1263
3 2 22 0 0 4224 0 21 19 0 0 4
773 1272
847 1272
847 1254
864 1254
3 1 23 0 0 8320 0 22 19 0 0 5
770 1202
770 1240
857 1240
857 1245
863 1245
1 0 11 0 0 0 0 22 0 0 100 2
725 1193
610 1193
2 0 10 0 0 0 0 22 0 0 110 2
725 1211
543 1211
1 0 10 0 0 0 0 21 0 0 110 2
728 1263
543 1263
0 2 9 0 0 0 0 0 21 111 0 3
505 1292
728 1292
728 1281
0 1 11 0 0 0 0 0 24 100 0 4
610 1087
711 1087
711 1080
721 1080
0 1 11 0 0 0 0 0 20 100 0 3
610 1340
610 1342
729 1342
2 0 9 0 0 0 0 20 0 0 111 2
729 1360
505 1360
0 1 9 0 0 0 0 0 23 111 0 4
505 1018
797 1018
797 1059
840 1059
2 3 24 0 0 4224 0 23 24 0 0 3
840 1077
770 1077
770 1089
2 0 10 0 0 0 0 24 0 0 110 2
721 1098
543 1098
5 2 25 0 0 8320 0 26 25 0 0 4
1016 746
1022 746
1022 684
1061 684
5 1 26 0 0 16512 0 27 25 0 0 6
1026 550
1030 550
1030 607
1029 607
1029 666
1061 666
3 0 27 0 0 4096 0 39 0 0 105 2
268 515
67 515
3 0 28 0 0 8192 0 28 0 0 66 3
663 777
663 778
661 778
3 0 29 0 0 8192 0 29 0 0 76 3
654 927
654 926
651 926
1 0 30 0 0 4096 0 36 0 0 109 2
271 733
156 733
1 0 30 0 0 4096 0 38 0 0 109 2
273 565
156 565
1 0 31 0 0 4096 0 39 0 0 104 2
268 497
221 497
2 0 32 0 0 4096 0 39 0 0 107 2
268 506
132 506
1 0 30 0 0 0 0 40 0 0 109 3
221 386
221 368
156 368
1 3 33 0 0 4224 0 51 52 0 0 4
700 500
664 500
664 499
656 499
0 2 10 0 0 0 0 0 52 110 0 2
543 508
611 508
0 1 9 0 0 0 0 0 52 111 0 2
505 490
611 490
2 4 34 0 0 12416 0 51 39 0 0 6
700 518
652 518
652 532
321 532
321 506
313 506
3 1 35 0 0 8320 0 51 27 0 0 5
745 509
745 510
914 510
914 537
976 537
3 1 36 0 0 4224 0 48 50 0 0 4
659 599
697 599
697 598
710 598
4 2 37 0 0 4224 0 38 50 0 0 4
318 574
702 574
702 616
710 616
3 2 38 0 0 4224 0 50 27 0 0 4
755 607
928 607
928 546
976 546
3 1 39 0 0 4224 0 49 47 0 0 2
657 699
723 699
0 2 10 0 0 0 0 0 49 110 0 2
543 708
611 708
0 1 9 0 0 0 0 0 49 111 0 2
505 690
611 690
0 2 10 0 0 0 0 0 48 110 0 2
543 608
608 608
0 1 9 0 0 0 0 0 48 111 0 2
505 590
608 590
4 2 40 0 0 4224 0 37 47 0 0 4
316 664
715 664
715 717
723 717
3 3 41 0 0 12416 0 27 47 0 0 6
976 555
935 555
935 633
781 633
781 708
768 708
1 0 28 0 0 4224 0 46 0 0 0 2
716 778
658 778
0 2 10 0 0 0 0 0 28 110 0 4
543 787
558 787
558 786
611 786
0 1 9 0 0 0 0 0 28 111 0 4
505 769
520 769
520 768
611 768
4 2 42 0 0 4224 0 36 46 0 0 4
316 742
703 742
703 796
716 796
4 3 43 0 0 8320 0 27 46 0 0 6
976 564
943 564
943 717
790 717
790 787
761 787
3 1 44 0 0 4224 0 45 44 0 0 2
648 852
713 852
0 2 9 0 0 0 0 0 45 111 0 2
505 861
599 861
0 1 10 0 0 0 0 0 45 110 0 2
543 843
599 843
4 2 45 0 0 4224 0 35 44 0 0 6
317 832
594 832
594 882
705 882
705 870
713 870
1 3 46 0 0 4224 0 26 44 0 0 4
966 733
802 733
802 861
758 861
0 1 29 0 0 4224 0 0 43 0 0 2
648 926
709 926
0 2 9 0 0 0 0 0 29 111 0 3
505 935
599 935
599 936
0 1 10 0 0 0 0 0 29 110 0 3
543 917
599 917
599 918
4 2 47 0 0 4224 0 34 43 0 0 6
307 909
594 909
594 956
701 956
701 944
709 944
3 2 48 0 0 8320 0 43 26 0 0 4
754 935
881 935
881 742
966 742
0 1 49 0 0 4096 0 0 42 106 0 3
39 378
67 378
67 381
0 1 50 0 0 4096 0 0 41 108 0 3
93 373
132 373
132 383
0 3 27 0 0 4096 0 0 38 105 0 2
67 583
273 583
0 2 32 0 0 4096 0 0 38 107 0 2
132 574
273 574
0 3 27 0 0 0 0 0 37 105 0 2
67 673
271 673
0 2 50 0 0 4096 0 0 37 108 0 2
93 664
271 664
0 3 27 0 0 0 0 0 36 105 0 2
67 751
271 751
0 2 50 0 0 0 0 0 36 108 0 2
93 742
271 742
0 3 49 0 0 4096 0 0 35 106 0 2
39 841
272 841
0 2 32 0 0 0 0 0 35 107 0 2
132 832
272 832
0 3 49 0 0 0 0 0 34 106 0 2
39 918
262 918
0 2 32 0 0 0 0 0 34 107 0 2
132 909
262 909
0 1 30 0 0 0 0 0 34 109 0 2
177 900
262 900
0 3 49 0 0 0 0 0 33 106 0 2
39 1131
258 1131
0 2 50 0 0 0 0 0 33 108 0 2
93 1122
258 1122
0 3 49 0 0 0 0 0 32 106 0 2
39 1256
259 1256
0 2 50 0 0 0 0 0 32 108 0 2
93 1247
259 1247
0 1 30 0 0 0 0 0 32 109 0 2
177 1238
259 1238
3 1 51 0 0 8320 0 25 31 0 0 4
1107 675
1107 674
1315 674
1315 649
1 0 11 0 0 12416 0 1 0 0 0 4
611 1053
611 1087
610 1087
610 1822
0 0 31 0 0 4096 0 0 0 102 0 2
221 1113
221 1402
1 0 31 0 0 8320 0 33 0 0 103 3
258 1113
221 1113
221 823
1 0 31 0 0 0 0 35 0 0 104 3
272 823
221 823
221 655
1 2 31 0 0 0 0 37 40 0 0 3
271 655
221 655
221 422
2 0 27 0 0 4224 0 42 0 0 0 2
67 417
67 1412
1 0 49 0 0 4224 0 4 0 0 0 2
39 359
39 1410
2 0 32 0 0 4224 0 41 0 0 0 2
132 419
132 1406
1 0 50 0 0 4224 0 3 0 0 0 2
93 361
93 1410
1 0 30 0 0 12416 0 2 0 0 0 4
156 359
156 738
177 738
177 1436
1 0 10 0 0 4224 0 5 0 0 0 2
543 476
543 1821
1 0 9 0 0 4224 0 6 0 0 0 2
505 476
505 1818
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
659 1465 736 1489
670 1474 724 1490
9 SUBTRADOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
682 990 747 1014
693 999 735 1015
7 SOMADOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
750 1165 785 1189
761 1174 773 1190
2 bc
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
735 1227 770 1251
746 1236 758 1252
2 ab
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
739 1303 774 1327
750 1312 762 1328
2 ac
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
493 390 578 405
507 401 563 412
8 ENTRADAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
49 266 141 281
63 277 126 288
9 CONTROLES
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
681 449 818 464
696 459 802 470
15 FUN�OES LOGICAS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
24 247 127 271
36 256 114 272
13 Decodificador
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
