CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 120 1 120 9
88 78 1856 788
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
46 800 1814 962
160432146 0
0
6 Title:
5 Name:
0
0
0
33
13 Logic Switch~
5 260 174 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-8 -22 6 -14
2 A3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 369 173 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-8 -22 6 -14
2 A2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 468 176 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-8 -22 6 -14
2 A1
-7 -30 7 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 569 172 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-8 -22 6 -14
2 A0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 177 439 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 ES
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 118 520 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 CLR
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 0 0 -2 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 170 239 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
5 CARGA
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9914 0 0
0
0
9 Inverter~
13 311 213 0 2 22
0 10 14
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
3747 0 0
0
0
9 Inverter~
13 419 211 0 2 22
0 11 15
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
3549 0 0
0
0
9 Inverter~
13 519 213 0 2 22
0 12 16
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
7931 0 0
0
0
9 Inverter~
13 617 209 0 2 22
0 13 18
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U6A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
9325 0 0
0
0
10 2-In NAND~
219 557 291 0 3 22
0 13 17 6
0
0 0 624 270
6 74LS00
-14 -24 28 -16
3 U5D
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
8903 0 0
0
0
10 2-In NAND~
219 609 292 0 3 22
0 18 17 2
0
0 0 624 270
6 74LS00
-14 -24 28 -16
3 U5C
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
3834 0 0
0
0
10 2-In NAND~
219 458 291 0 3 22
0 12 17 7
0
0 0 624 270
6 74LS00
-14 -24 28 -16
3 U5B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
3363 0 0
0
0
10 2-In NAND~
219 510 292 0 3 22
0 16 17 3
0
0 0 624 270
6 74LS00
-14 -24 28 -16
3 U5A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
7668 0 0
0
0
10 2-In NAND~
219 358 290 0 3 22
0 11 17 8
0
0 0 624 270
6 74LS00
-14 -24 28 -16
3 U4D
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
4718 0 0
0
0
10 2-In NAND~
219 410 291 0 3 22
0 15 17 4
0
0 0 624 270
6 74LS00
-14 -24 28 -16
3 U4C
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3874 0 0
0
0
10 2-In NAND~
219 301 297 0 3 22
0 14 17 5
0
0 0 624 270
6 74LS00
-14 -24 28 -16
3 U4B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6671 0 0
0
0
10 2-In NAND~
219 249 296 0 3 22
0 10 17 9
0
0 0 624 270
6 74LS00
-14 -24 28 -16
3 U4A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3789 0 0
0
0
14 Logic Display~
6 640 341 0 1 2
10 20
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 535 339 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3750 0 0
0
0
14 Logic Display~
6 429 338 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8778 0 0
0
0
5 SCOPE
12 647 406 0 1 11
0 20
0
0 0 57584 270
2 Q4
-8 -4 6 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
538 0 0
0
0
5 SCOPE
12 544 407 0 1 11
0 21
0
0 0 57584 270
2 Q3
-8 -4 6 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
6843 0 0
0
0
5 SCOPE
12 436 407 0 1 11
0 22
0
0 0 57584 270
2 Q2
-8 -4 6 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
3136 0 0
0
0
5 SCOPE
12 341 399 0 1 11
0 19
0
0 0 57584 270
2 Q1
-8 -4 6 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
5950 0 0
0
0
5 7474~
219 581 475 0 6 22
0 6 21 23 2 26 20
0
0 0 4720 0
6 74LS74
0 -60 42 -52
3 U1B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
65 0 0 512 2 2 3 0
1 U
5670 0 0
0
0
5 7474~
219 482 476 0 6 22
0 7 22 23 3 27 21
0
0 0 4720 0
6 74LS74
0 -60 42 -52
3 U1A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
65 0 0 512 2 1 3 0
1 U
6828 0 0
0
0
5 7474~
219 368 474 0 6 22
0 8 19 23 4 28 22
0
0 0 4720 0
6 74LS74
0 -60 42 -52
3 U3B
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 10 12 11 13 8 9 4 2 3
1 6 5 10 12 11 13 8 9 0
65 0 0 512 2 2 2 0
1 U
6735 0 0
0
0
5 7474~
219 251 476 0 6 22
0 9 24 23 5 29 19
0
0 0 4720 0
6 74LS74
0 -60 42 -52
3 U3A
22 -61 43 -53
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 4 2 3 1 6 5 4 2 3
1 6 5 10 12 11 13 8 9 0
65 0 0 512 2 1 2 0
1 U
8365 0 0
0
0
5 SCOPE
12 177 477 0 1 11
0 23
0
0 0 57584 270
2 CK
-7 -4 7 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
0
4132 0 0
0
0
7 Pulser~
4 109 463 0 10 12
0 30 31 23 32 0 0 5 5 5
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4551 0 0
0
0
14 Logic Display~
6 334 335 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3635 0 0
0
0
51
3 4 2 0 0 8336 0 13 27 0 0 4
610 318
621 318
621 487
581 487
3 4 3 0 0 4224 0 15 28 0 0 6
511 318
511 409
453 409
453 496
482 496
482 488
3 4 4 0 0 4224 0 17 29 0 0 4
411 317
411 494
368 494
368 486
3 4 5 0 0 4224 0 18 30 0 0 4
302 323
302 496
251 496
251 488
3 1 6 0 0 4224 0 12 27 0 0 4
558 317
558 404
581 404
581 412
3 1 7 0 0 4224 0 14 28 0 0 4
459 317
459 405
482 405
482 413
1 3 8 0 0 4224 0 29 16 0 0 3
368 411
368 316
359 316
3 1 9 0 0 8320 0 19 30 0 0 3
250 322
251 322
251 413
1 0 10 0 0 4096 0 1 0 0 13 2
260 186
261 186
1 0 11 0 0 4096 0 2 0 0 16 2
369 185
369 184
1 0 12 0 0 4096 0 3 0 0 21 2
468 188
469 186
1 0 13 0 0 4096 0 4 0 0 31 2
569 184
569 182
1 1 10 0 0 12416 0 8 19 0 0 5
314 195
314 186
261 186
261 271
259 271
2 0 14 0 0 4096 0 8 0 0 15 2
314 231
313 231
1 0 14 0 0 8320 0 18 0 0 0 3
311 272
313 272
313 228
1 1 11 0 0 12416 0 9 16 0 0 5
422 193
422 184
369 184
369 265
368 265
2 0 15 0 0 4096 0 9 0 0 18 2
422 229
421 229
1 0 15 0 0 8320 0 17 0 0 0 3
420 266
421 266
421 226
1 0 16 0 0 4096 0 15 0 0 23 2
520 267
521 267
1 0 12 0 0 0 0 14 0 0 21 2
468 266
469 266
1 1 12 0 0 12416 0 10 0 0 0 4
522 195
522 186
469 186
469 270
2 0 16 0 0 0 0 10 0 0 23 2
522 231
521 231
1 0 16 0 0 4224 0 0 0 0 0 2
521 271
521 228
2 0 17 0 0 4096 0 16 0 0 34 4
350 265
350 242
349 242
349 239
2 0 17 0 0 4096 0 19 0 0 34 2
241 271
241 239
0 2 17 0 0 4096 0 0 18 34 0 3
296 239
296 272
293 272
2 0 17 0 0 0 0 17 0 0 34 2
402 266
402 239
2 0 17 0 0 0 0 14 0 0 34 2
450 266
450 239
2 0 17 0 0 0 0 15 0 0 34 2
502 267
502 239
2 0 17 0 0 0 0 12 0 0 34 2
549 266
549 239
1 1 13 0 0 12416 0 11 12 0 0 4
620 191
620 182
567 182
567 266
2 0 18 0 0 4096 0 11 0 0 33 2
620 227
619 227
1 0 18 0 0 4224 0 13 0 0 0 2
619 267
619 224
1 2 17 0 0 4224 0 7 13 0 0 3
182 239
601 239
601 267
0 1 19 0 0 4224 0 0 33 51 0 3
335 438
335 353
334 353
1 0 20 0 0 4096 0 23 0 0 44 2
638 409
640 409
1 0 21 0 0 4096 0 24 0 0 45 2
535 410
536 410
1 0 22 0 0 4096 0 25 0 0 46 2
427 410
428 410
1 0 19 0 0 0 0 26 0 0 35 4
332 402
321 402
321 405
335 405
1 0 23 0 0 0 0 31 0 0 43 2
168 480
168 480
3 0 23 0 0 8192 0 28 0 0 43 3
458 458
447 458
447 507
3 0 23 0 0 8192 0 29 0 0 43 3
344 456
332 456
332 507
0 3 23 0 0 8320 0 0 27 47 0 4
168 454
168 507
557 507
557 457
6 1 20 0 0 8320 0 27 20 0 0 3
605 439
640 439
640 359
0 1 21 0 0 4224 0 0 21 49 0 3
536 439
536 357
535 357
0 1 22 0 0 4224 0 0 22 50 0 3
428 440
428 356
429 356
3 3 23 0 0 0 0 32 30 0 0 4
133 454
219 454
219 458
227 458
2 1 24 0 0 4224 0 30 5 0 0 3
227 440
189 440
189 439
6 2 21 0 0 0 0 28 27 0 0 3
506 440
506 439
557 439
6 2 22 0 0 0 0 29 28 0 0 3
392 438
392 440
458 440
6 2 19 0 0 0 0 30 29 0 0 3
275 440
275 438
344 438
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
