CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
617 143 1863 1128
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
51 C:\Users\guipa\OneDrive\�rea de Trabalho\cm\BOM.DAT
0 7
0 4 0.500000 0.500000
785 239 898 336
42991634 0
0
6 Title:
5 Name:
0
0
0
34
13 Logic Switch~
5 152 345 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4874 0 0
2
5.89923e-315 0
0
13 Logic Switch~
5 256 644 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
886 0 0
2
5.89923e-315 5.30499e-315
0
13 Logic Switch~
5 259 678 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3181 0 0
2
5.89923e-315 5.26354e-315
0
13 Logic Switch~
5 256 716 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5363 0 0
2
5.89923e-315 0
0
13 Logic Switch~
5 257 120 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5407 0 0
2
5.89923e-315 0
0
13 Logic Switch~
5 260 82 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4378 0 0
2
5.89923e-315 0
0
13 Logic Switch~
5 257 48 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6531 0 0
2
5.89923e-315 0
0
5 4081~
219 830 707 0 3 22
0 8 7 11
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U11D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
9150 0 0
2
5.89923e-315 0
0
5 4081~
219 831 649 0 3 22
0 9 7 12
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U11C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
4532 0 0
2
5.89923e-315 0
0
5 4081~
219 826 599 0 3 22
0 10 7 13
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U11B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
3472 0 0
2
5.89923e-315 0
0
5 4073~
219 399 736 0 4 22
0 16 15 14 7
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
8894 0 0
2
5.89923e-315 0
0
5 4071~
219 743 524 0 3 22
0 18 19 10
0
0 0 624 270
4 4071
-7 -24 21 -16
3 U9C
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
9568 0 0
2
5.89923e-315 0
0
5 4071~
219 583 522 0 3 22
0 20 21 9
0
0 0 624 270
4 4071
-7 -24 21 -16
3 U9B
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
9334 0 0
2
5.89923e-315 0
0
5 4071~
219 434 520 0 3 22
0 26 25 8
0
0 0 624 270
4 4071
-7 -24 21 -16
3 U9A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3276 0 0
2
5.89923e-315 0
0
5 4049~
219 250 263 0 2 22
0 2 3
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U12F
-8 -21 20 -13
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 6 0
1 U
3252 0 0
2
5.89923e-315 0
0
14 Logic Display~
6 893 695 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
530 0 0
2
5.89923e-315 0
0
14 Logic Display~
6 895 648 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5772 0 0
2
5.89923e-315 0
0
14 Logic Display~
6 893 596 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4918 0 0
2
5.89923e-315 0
0
5 4049~
219 362 617 0 2 22
0 15 17
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U12A
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 6 0
1 U
6443 0 0
2
5.89923e-315 0
0
5 4081~
219 787 427 0 3 22
0 24 2 19
0
0 0 624 270
4 4081
-7 -24 21 -16
4 U11A
13 -4 41 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
4904 0 0
2
5.89923e-315 0
0
5 4081~
219 809 268 0 3 22
0 29 3 18
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U8D
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
5677 0 0
2
5.89923e-315 0
0
5 4081~
219 369 527 0 3 22
0 16 17 6
0
0 0 624 90
4 4081
-7 -24 21 -16
3 U8C
16 -5 37 3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
4454 0 0
2
5.89923e-315 0
0
5 4081~
219 625 428 0 3 22
0 23 2 21
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U8B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
5604 0 0
2
5.89923e-315 0
0
5 4081~
219 463 427 0 3 22
0 22 2 25
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U8A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3284 0 0
2
5.89923e-315 0
0
5 4081~
219 653 269 0 3 22
0 27 3 20
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U7D
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
9222 0 0
2
5.89923e-315 0
0
5 4081~
219 496 273 0 3 22
0 28 3 26
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U7C
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
9672 0 0
2
5.89923e-315 0
0
5 4081~
219 323 389 0 3 22
0 2 6 4
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
996 0 0
2
5.89923e-315 0
0
5 4081~
219 317 240 0 3 22
0 6 3 5
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
8631 0 0
2
5.89923e-315 0
0
12 D Flip-Flop~
219 714 379 0 4 9
0 32 4 33 24
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U6
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9515 0 0
2
5.89923e-315 0
0
12 D Flip-Flop~
219 564 380 0 4 9
0 31 4 34 23
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U5
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7604 0 0
2
5.89923e-315 0
0
12 D Flip-Flop~
219 417 379 0 4 9
0 30 4 35 22
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U4
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9545 0 0
2
5.89923e-315 0
0
12 D Flip-Flop~
219 717 235 0 4 9
0 32 5 36 29
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U3
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8952 0 0
2
5.89923e-315 0
0
12 D Flip-Flop~
219 564 236 0 4 9
0 31 5 37 27
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U2
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8283 0 0
2
5.89923e-315 0
0
12 D Flip-Flop~
219 416 239 0 4 9
0 30 5 38 28
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4938 0 0
2
5.89923e-315 0
0
51
0 0 2 0 0 4096 0 0 0 9 3 2
164 351
235 351
2 2 3 0 0 4096 0 28 15 0 0 4
293 249
279 249
279 263
271 263
1 1 2 0 0 4096 0 15 27 0 0 3
235 263
235 380
299 380
2 2 3 0 0 8192 0 25 21 0 0 3
642 247
642 246
798 246
2 2 3 0 0 8192 0 26 25 0 0 3
485 251
485 247
642 247
2 2 3 0 0 4224 0 15 26 0 0 4
271 263
470 263
470 251
485 251
0 2 2 0 0 8192 0 0 20 8 0 4
612 398
612 392
776 392
776 405
2 2 2 0 0 0 0 24 23 0 0 4
452 405
452 398
614 398
614 406
1 2 2 0 0 8320 0 1 24 0 0 3
164 345
164 405
452 405
0 0 4 0 0 8192 0 0 0 12 13 3
539 389
539 385
686 385
3 0 4 0 0 0 0 27 0 0 12 2
344 389
372 389
2 2 4 0 0 12416 0 31 30 0 0 5
393 361
372 361
372 389
540 389
540 362
2 0 4 0 0 0 0 29 0 0 0 3
690 361
686 361
686 389
0 2 5 0 0 4224 0 0 32 15 0 4
531 240
685 240
685 217
693 217
0 2 5 0 0 0 0 0 33 16 0 4
384 240
532 240
532 218
540 218
3 2 5 0 0 0 0 28 34 0 0 4
338 240
384 240
384 221
392 221
1 0 6 0 0 8320 0 28 0 0 18 4
293 231
205 231
205 496
295 496
2 3 6 0 0 0 0 27 22 0 0 5
299 398
295 398
295 496
368 496
368 503
0 2 7 0 0 4096 0 0 10 21 0 3
698 736
698 608
802 608
0 2 7 0 0 0 0 0 9 21 0 3
752 736
752 658
807 658
4 2 7 0 0 4224 0 11 8 0 0 4
420 736
798 736
798 716
806 716
3 1 8 0 0 8320 0 14 8 0 0 3
437 550
437 698
806 698
1 3 9 0 0 4224 0 9 13 0 0 3
807 640
586 640
586 552
1 3 10 0 0 4224 0 10 12 0 0 3
802 590
746 590
746 554
3 1 11 0 0 4224 0 8 16 0 0 5
851 707
881 707
881 721
893 721
893 713
3 1 12 0 0 4224 0 9 17 0 0 5
852 649
883 649
883 674
895 674
895 666
3 1 13 0 0 4224 0 10 18 0 0 5
847 599
881 599
881 622
893 622
893 614
1 3 14 0 0 8320 0 4 11 0 0 3
268 716
268 745
375 745
0 2 15 0 0 8192 0 0 11 31 0 3
298 678
298 736
375 736
0 1 16 0 0 4224 0 0 11 33 0 3
325 559
325 727
375 727
1 1 15 0 0 4224 0 3 19 0 0 3
271 678
365 678
365 635
2 2 17 0 0 4224 0 19 22 0 0 4
365 599
365 562
377 562
377 548
1 1 16 0 0 0 0 2 22 0 0 4
268 644
268 559
359 559
359 548
1 3 18 0 0 12416 0 12 21 0 0 4
755 508
755 498
807 498
807 291
2 3 19 0 0 8320 0 12 20 0 0 4
737 508
737 486
785 486
785 450
1 3 20 0 0 8320 0 13 25 0 0 3
595 506
651 506
651 292
3 2 21 0 0 8320 0 23 13 0 0 4
623 451
623 492
577 492
577 506
1 4 22 0 0 4224 0 24 31 0 0 3
470 405
470 343
441 343
1 4 23 0 0 4224 0 23 30 0 0 3
632 406
632 344
588 344
1 4 24 0 0 4224 0 20 29 0 0 3
794 405
794 343
738 343
3 2 25 0 0 12416 0 24 14 0 0 4
461 450
461 470
428 470
428 504
1 3 26 0 0 12416 0 14 26 0 0 4
446 504
446 480
494 480
494 296
1 4 27 0 0 8320 0 25 33 0 0 3
660 247
660 200
588 200
1 4 28 0 0 8320 0 26 34 0 0 3
503 251
503 203
440 203
4 1 29 0 0 4224 0 32 21 0 0 3
741 199
816 199
816 246
0 1 30 0 0 8192 0 0 34 47 0 4
380 212
386 212
386 203
392 203
1 1 30 0 0 8320 0 5 31 0 0 4
269 120
380 120
380 343
393 343
0 1 31 0 0 8192 0 0 33 49 0 3
527 212
527 200
540 200
1 1 31 0 0 8320 0 6 30 0 0 4
272 82
527 82
527 344
540 344
0 1 32 0 0 8192 0 0 32 51 0 3
677 211
677 199
693 199
1 1 32 0 0 4224 0 7 29 0 0 4
269 48
677 48
677 343
690 343
8
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
886 533 1019 562
896 541 1008 560
14 Sa�da de dados
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
202 700 239 729
212 708 228 727
2 OE
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
202 662 239 691
212 670 228 689
2 RD
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
203 629 240 658
213 637 229 656
2 CS
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 16
160 -5 309 24
170 3 298 22
16 Entrada de dados
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 11
24 324 133 353
34 332 122 351
11 Controlador
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
822 342 915 371
832 350 904 369
9 Palavra 2
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
821 206 914 235
831 214 903 233
9 Palavra 1
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
