CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 120 3 120 9
88 78 1856 788
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
88 78 1856 788
143654930 0
0
6 Title:
5 Name:
0
0
0
27
13 Logic Switch~
5 272 462 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -17 9 -9
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 336 253 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -17 9 -9
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 348 298 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -17 9 -9
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 351 407 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -17 9 -9
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
9 Inverter~
13 392 407 0 2 22
0 18 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U6A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
5394 0 0
0
0
9 2-In AND~
219 958 321 0 3 22
0 17 3 12
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
7734 0 0
0
0
9 2-In AND~
219 959 369 0 3 22
0 6 18 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
9914 0 0
0
0
8 2-In OR~
219 1009 342 0 3 22
0 12 11 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
3747 0 0
0
0
9 2-In AND~
219 757 321 0 3 22
0 17 4 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
3549 0 0
0
0
9 2-In AND~
219 758 369 0 3 22
0 7 18 13
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
7931 0 0
0
0
8 2-In OR~
219 808 342 0 3 22
0 14 13 21
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9325 0 0
0
0
8 2-In OR~
219 594 338 0 3 22
0 16 15 9
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
8903 0 0
0
0
9 2-In AND~
219 544 365 0 3 22
0 20 18 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3834 0 0
0
0
9 2-In AND~
219 543 317 0 3 22
0 17 5 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3363 0 0
0
0
14 Logic Display~
6 929 187 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7668 0 0
0
0
14 Logic Display~
6 810 185 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
14 Logic Display~
6 664 184 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3874 0 0
0
0
14 Logic Display~
6 519 187 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6671 0 0
0
0
14 Logic Display~
6 785 483 0 1 2
10 24
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L4
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3789 0 0
0
0
14 Logic Display~
6 917 495 0 1 2
10 25
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 654 493 0 1 2
10 26
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3750 0 0
0
0
14 Logic Display~
6 507 494 0 1 2
10 27
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
8778 0 0
0
0
7 Pulser~
4 251 352 0 10 12
0 28 29 23 30 0 0 5 5 1
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
538 0 0
0
0
6 74112~
219 1100 368 0 7 32
0 22 8 10 8 19 31 2
0
0 0 4720 0
6 74LS76
0 -60 42 -52
3 U2B
22 -61 43 -53
0
15 DVCC=5;DGND=13;
72 %D [%5bi %13bi %1i %2i %3i %4i %5i][%5bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 9 6 12 8 10 11 2 4
1 16 3 14 15 7 9 6 12 8
10 11 0
65 0 0 512 2 2 2 0
1 U
6843 0 0
0
0
6 74112~
219 882 369 0 7 32
0 22 8 21 8 19 6 3
0
0 0 4720 0
6 74LS76
0 -60 42 -52
3 U2A
22 -61 43 -53
0
15 DVCC=5;DGND=13;
72 %D [%5bi %13bi %1i %2i %3i %4i %5i][%5bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 2 4 1 16 3 14 15 2 4
1 16 3 14 15 7 9 6 12 8
10 11 0
65 0 0 0 2 1 2 0
1 U
3136 0 0
0
0
6 74112~
219 680 366 0 7 32
0 22 8 9 8 19 7 4
0
0 0 4720 0
6 74LS76
0 -60 42 -52
3 U1B
22 -61 43 -53
0
15 DVCC=5;DGND=13;
72 %D [%5bi %13bi %1i %2i %3i %4i %5i][%5bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 9 6 12 8 10 11 2 4
1 16 3 14 15 7 9 6 12 8
10 11 0
65 0 0 0 2 2 1 0
1 U
5950 0 0
0
0
6 74112~
219 473 375 0 7 32
0 22 8 23 8 19 20 5
0
0 0 4720 0
6 74LS76
0 -60 42 -52
3 U1A
22 -61 43 -53
0
15 DVCC=5;DGND=13;
72 %D [%5bi %13bi %1i %2i %3i %4i %5i][%5bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 2 4 1 16 3 14 15 2 4
1 16 3 14 15 7 9 6 12 8
10 11 1270830282
65 0 0 0 2 1 1 0
1 U
5670 0 0
0
0
44
7 1 2 0 0 8320 0 24 15 0 0 3
1124 332
1124 205
929 205
0 1 3 0 0 12416 0 0 16 6 0 6
914 333
914 385
790 385
790 211
810 211
810 203
0 1 4 0 0 12416 0 0 17 7 0 6
710 330
710 382
645 382
645 210
664 210
664 202
0 1 5 0 0 12416 0 0 18 35 0 6
502 339
502 391
515 391
515 213
519 213
519 205
1 6 6 0 0 4224 0 7 25 0 0 4
935 360
920 360
920 351
912 351
2 7 3 0 0 0 0 6 25 0 0 4
934 330
920 330
920 333
906 333
7 2 4 0 0 0 0 26 9 0 0 2
704 330
733 330
6 1 7 0 0 4224 0 26 10 0 0 4
710 348
726 348
726 360
734 360
2 0 8 0 0 8192 0 26 0 0 12 3
656 330
646 330
646 298
2 0 8 0 0 8192 0 25 0 0 12 3
858 333
848 333
848 298
0 2 8 0 0 4096 0 0 27 12 0 3
435 298
435 339
449 339
1 2 8 0 0 4224 0 3 24 0 0 4
360 298
1062 298
1062 332
1076 332
4 2 8 0 0 0 0 26 26 0 0 4
656 348
642 348
642 330
656 330
4 2 8 0 0 0 0 25 25 0 0 4
858 351
846 351
846 333
858 333
4 2 8 0 0 0 0 24 24 0 0 4
1076 350
1062 350
1062 332
1076 332
3 3 9 0 0 4224 0 12 26 0 0 4
627 338
642 338
642 339
650 339
3 3 10 0 0 4224 0 8 24 0 0 4
1042 342
1062 342
1062 341
1070 341
2 3 11 0 0 8320 0 8 7 0 0 4
996 351
988 351
988 369
980 369
3 1 12 0 0 8320 0 6 8 0 0 4
979 321
988 321
988 333
996 333
2 3 13 0 0 8320 0 11 10 0 0 4
795 351
787 351
787 369
779 369
1 3 14 0 0 8320 0 11 9 0 0 4
795 333
786 333
786 321
778 321
2 3 15 0 0 8320 0 12 13 0 0 4
581 347
573 347
573 365
565 365
1 3 16 0 0 8320 0 12 14 0 0 4
581 329
572 329
572 317
564 317
1 0 17 0 0 8192 0 14 0 0 32 3
519 308
508 308
508 407
1 0 17 0 0 0 0 9 0 0 32 3
733 312
714 312
714 407
2 0 18 0 0 8192 0 10 0 0 33 3
734 378
730 378
730 451
2 0 18 0 0 8192 0 13 0 0 33 3
520 374
516 374
516 451
5 0 19 0 0 4096 0 25 0 0 31 2
882 381
882 463
5 0 19 0 0 4096 0 26 0 0 31 2
680 378
680 463
5 0 19 0 0 0 0 27 0 0 31 2
473 387
473 463
5 1 19 0 0 8320 0 24 1 0 0 4
1100 380
1100 463
284 463
284 462
2 1 17 0 0 4224 0 5 6 0 0 4
413 407
926 407
926 312
934 312
0 2 18 0 0 8320 0 0 7 44 0 4
370 407
370 451
935 451
935 378
6 1 20 0 0 4224 0 27 13 0 0 4
503 357
512 357
512 356
520 356
7 2 5 0 0 0 0 27 14 0 0 4
497 339
511 339
511 326
519 326
3 3 21 0 0 4224 0 25 11 0 0 2
852 342
841 342
1 0 22 0 0 0 0 2 0 0 41 2
348 253
348 253
1 0 22 0 0 8192 0 25 0 0 41 4
882 306
882 268
756 268
756 253
1 0 22 0 0 0 0 26 0 0 41 4
680 303
680 268
623 268
623 253
1 0 22 0 0 0 0 27 0 0 41 2
473 312
473 253
1 0 22 0 0 8320 0 24 0 0 0 3
1100 305
1100 253
344 253
3 3 23 0 0 4224 0 23 27 0 0 4
275 343
435 343
435 348
443 348
4 2 8 0 0 0 0 27 27 0 0 4
449 357
432 357
432 339
449 339
1 1 18 0 0 128 0 4 5 0 0 2
363 407
377 407
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
