CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 4 90 10
189 83 1534 801
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
357 179 470 276
42991634 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 321 267 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7290 0 0
2
5.89924e-315 0
0
13 Logic Switch~
5 179 694 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3576 0 0
2
43847.9 0
0
5 4081~
219 519 924 0 3 22
0 5 4 3
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U2C
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
7787 0 0
2
5.89924e-315 0
0
5 4081~
219 676 226 0 3 22
0 6 7 9
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
7379 0 0
2
43847.9 1
0
5 4081~
219 510 229 0 3 22
0 6 11 10
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
5233 0 0
2
43847.9 2
0
6 JK RN~
219 728 339 0 6 22
0 9 3 6 12 11 8
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 1 4 0
1 U
4421 0 0
2
43847.9 3
0
6 JK RN~
219 588 341 0 6 22
0 10 3 6 12 20 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 3 0
1 U
3157 0 0
2
43847.9 4
0
6 JK RN~
219 444 337 0 6 22
0 12 3 12 12 21 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 3 0
1 U
7411 0 0
2
43847.9 5
0
12 Hex Display~
7 961 212 0 16 19
10 6 7 8 22 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
8362 0 0
2
5.89924e-315 5.30499e-315
0
12 Hex Display~
7 1014 210 0 16 19
10 4 13 14 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3199 0 0
2
43847.9 6
0
5 4073~
219 647 580 0 4 22
0 4 13 14 15
0
0 0 624 270
4 4073
-7 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
4127 0 0
2
43847.9 7
0
7 Pulser~
4 111 757 0 10 12
0 23 24 19 25 0 0 10 10 11
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7649 0 0
2
43847.9 8
0
6 74112~
219 775 783 0 7 32
0 2 15 19 4 2 16 5
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 3 0
1 U
5225 0 0
2
43847.9 9
0
6 74112~
219 615 784 0 7 32
0 2 17 19 26 2 27 14
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
4702 0 0
2
43847.9 10
0
6 74112~
219 444 793 0 7 32
0 2 18 19 4 2 28 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
60 0 0
2
43847.9 11
0
6 74112~
219 277 791 0 7 32
0 2 2 19 2 2 29 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
5704 0 0
2
43847.9 12
0
5 4081~
219 500 585 0 3 22
0 4 13 17
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U1B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
4208 0 0
2
43847.9 13
0
5 4081~
219 364 586 0 3 22
0 16 4 18
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U1A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3666 0 0
2
43847.9 14
0
56
0 0 2 0 0 8192 0 0 0 8 9 3
615 991
628 991
628 1005
0 0 2 0 0 8192 0 0 0 9 52 3
278 1005
212 1005
212 694
0 0 3 0 0 8192 0 0 0 6 4 3
351 336
351 329
343 329
3 2 3 0 0 12416 0 3 8 0 0 5
517 947
517 1044
71 1044
71 329
413 329
0 2 4 0 0 4096 0 0 3 31 0 6
305 755
305 954
497 954
497 894
508 894
508 902
0 0 3 0 0 0 0 0 0 12 0 2
351 344
351 329
5 0 2 0 0 0 0 15 0 0 9 2
444 805
444 1005
5 0 2 0 0 0 0 14 0 0 0 4
615 796
615 1000
616 1000
616 1005
5 5 2 0 0 8192 0 13 16 0 0 4
775 795
775 1005
277 1005
277 803
1 0 5 0 0 16384 0 3 0 0 11 6
526 902
526 894
537 894
537 954
808 954
808 747
7 4 5 0 0 8320 0 13 10 0 0 3
799 747
1005 747
1005 234
0 0 3 0 0 0 0 0 0 57 13 3
351 341
351 349
365 349
0 2 3 0 0 0 0 0 6 0 0 4
365 344
365 448
697 448
697 331
1 6 6 0 0 8320 0 9 8 0 0 5
970 236
970 297
491 297
491 320
468 320
2 0 7 0 0 8320 0 9 0 0 19 3
964 236
964 302
612 302
3 6 8 0 0 8320 0 9 6 0 0 3
958 236
958 322
752 322
3 1 9 0 0 4224 0 4 6 0 0 3
697 226
697 322
704 322
1 0 6 0 0 0 0 4 0 0 24 5
652 217
542 217
542 199
468 199
468 221
6 2 7 0 0 0 0 7 4 0 0 3
612 324
612 235
652 235
3 1 10 0 0 4224 0 5 7 0 0 3
531 229
531 324
564 324
2 5 11 0 0 8320 0 5 6 0 0 5
486 238
486 287
769 287
769 340
758 340
3 0 6 0 0 0 0 7 0 0 23 2
564 342
485 342
6 3 6 0 0 0 0 8 6 0 0 5
468 320
485 320
485 377
704 377
704 340
6 1 6 0 0 0 0 8 5 0 0 5
468 320
468 221
472 221
472 220
486 220
4 0 12 0 0 4096 0 8 0 0 27 4
444 368
444 383
448 383
448 391
4 0 12 0 0 4096 0 7 0 0 27 2
588 372
588 391
0 4 12 0 0 8320 0 0 6 28 0 4
409 344
409 391
728 391
728 370
0 3 12 0 0 0 0 0 8 29 0 5
409 326
409 344
409 344
409 338
420 338
1 1 12 0 0 0 0 1 8 0 0 6
333 267
409 267
409 326
409 326
409 320
420 320
2 0 3 0 0 0 0 7 0 0 13 3
557 333
554 333
554 448
1 0 4 0 0 8320 0 10 0 0 42 4
1023 234
1023 705
305 705
305 755
2 0 13 0 0 8320 0 10 0 0 40 4
1017 234
1017 710
472 710
472 757
3 7 14 0 0 4224 0 10 14 0 0 5
1011 234
1011 715
653 715
653 748
639 748
0 0 4 0 0 0 0 0 0 35 44 4
524 544
398 544
398 645
326 645
1 0 4 0 0 0 0 11 0 0 39 5
654 558
654 544
523 544
523 553
506 553
2 0 13 0 0 0 0 11 0 0 40 4
645 558
645 535
485 535
485 563
3 7 14 0 0 0 0 11 14 0 0 9
636 558
636 546
612 546
612 652
626 652
626 678
669 678
669 748
639 748
4 2 15 0 0 12416 0 11 13 0 0 6
645 603
645 655
718 655
718 743
751 743
751 747
0 1 4 0 0 0 0 0 17 44 0 5
326 624
430 624
430 553
507 553
507 563
2 7 13 0 0 0 0 17 15 0 0 4
489 563
477 563
477 757
468 757
1 6 16 0 0 8320 0 18 13 0 0 5
371 564
371 530
911 530
911 765
805 765
7 0 4 0 0 0 0 16 0 0 44 2
301 755
326 755
0 4 4 0 0 0 0 0 15 44 0 2
326 775
420 775
2 4 4 0 0 0 0 18 13 0 0 5
353 564
326 564
326 870
751 870
751 765
3 2 17 0 0 4224 0 17 14 0 0 3
498 608
498 748
591 748
3 2 18 0 0 4224 0 18 15 0 0 3
362 609
362 757
420 757
0 4 2 0 0 0 0 0 16 48 0 4
227 755
234 755
234 773
253 773
0 2 2 0 0 0 0 0 16 52 0 3
227 694
227 755
253 755
0 1 2 0 0 0 0 0 16 52 0 2
277 694
277 728
0 1 2 0 0 0 0 0 15 52 0 2
444 694
444 730
0 1 2 0 0 0 0 0 14 52 0 2
615 694
615 721
1 1 2 0 0 4224 0 2 13 0 0 3
191 694
775 694
775 720
3 0 19 0 0 8192 0 15 0 0 55 3
414 766
410 766
410 883
3 0 19 0 0 8192 0 14 0 0 55 3
585 757
577 757
577 883
0 3 19 0 0 8320 0 0 13 56 0 4
185 748
185 883
745 883
745 756
3 3 19 0 0 0 0 12 16 0 0 4
135 748
239 748
239 764
247 764
2
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 15
396 484 679 532
409 493 665 525
15 Circuito MOD-10
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
429 150 694 198
442 159 680 191
14 Circuito MOD-6
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
