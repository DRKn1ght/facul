CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 60 1 90 10
1983 189 3229 1149
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
2 4 0.500000 0.500000
2151 285 2264 382
9437202 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 321 267 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7145 0 0
2
5.89923e-315 0
0
13 Logic Switch~
5 179 694 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6215 0 0
2
43844.8 0
0
5 4011~
219 519 979 0 3 22
0 4 2 3
0
0 0 624 270
4 4011
-7 -24 21 -16
3 U5A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 6 0
1 U
664 0 0
2
5.89923e-315 0
0
5 4081~
219 676 226 0 3 22
0 5 6 8
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
9523 0 0
2
43844.8 1
0
5 4081~
219 510 229 0 3 22
0 5 10 9
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
7629 0 0
2
43844.8 2
0
6 JK RN~
219 728 339 0 6 22
0 8 3 5 11 10 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 1 4 0
1 U
5231 0 0
2
43844.8 3
0
6 JK RN~
219 588 341 0 6 22
0 9 3 5 11 20 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 3 0
1 U
360 0 0
2
43844.8 4
0
6 JK RN~
219 444 337 0 6 22
0 11 3 11 11 21 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 3 0
1 U
3318 0 0
2
43844.8 5
0
12 Hex Display~
7 961 212 0 16 19
10 5 6 7 22 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
8169 0 0
2
5.89923e-315 5.30499e-315
0
12 Hex Display~
7 1014 210 0 16 19
10 2 12 13 4 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3347 0 0
2
43844.8 6
0
5 4073~
219 647 580 0 4 22
0 2 12 13 14
0
0 0 624 270
4 4073
-7 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
9798 0 0
2
43844.8 7
0
7 Pulser~
4 111 757 0 10 12
0 23 24 19 25 0 0 10 10 11
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3254 0 0
2
43844.8 8
0
6 74112~
219 775 783 0 7 32
0 18 14 19 2 3 15 4
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 2 3 0
1 U
5152 0 0
2
43844.8 9
0
6 74112~
219 615 784 0 7 32
0 18 16 19 26 3 27 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
756 0 0
2
43844.8 10
0
6 74112~
219 444 793 0 7 32
0 18 17 19 2 3 28 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3391 0 0
2
43844.8 11
0
6 74112~
219 277 791 0 7 32
0 18 18 19 18 3 29 2
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
986 0 0
2
43844.8 12
0
5 4081~
219 500 585 0 3 22
0 2 12 16
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U1B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
9485 0 0
2
43844.8 13
0
5 4081~
219 364 586 0 3 22
0 15 2 17
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U1A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3897 0 0
2
43844.8 14
0
54
0 2 2 0 0 8192 0 0 3 29 0 3
305 755
305 954
511 954
0 0 3 0 0 4096 0 0 0 10 3 2
351 344
351 329
3 2 3 0 0 12416 0 3 8 0 0 5
520 1005
520 1027
64 1027
64 329
413 329
5 0 3 0 0 0 0 15 0 0 7 2
444 805
444 1005
5 0 3 0 0 0 0 14 0 0 6 4
615 796
615 1000
616 1000
616 1005
3 5 3 0 0 0 0 3 13 0 0 3
520 1005
775 1005
775 795
3 5 3 0 0 0 0 3 16 0 0 3
520 1005
277 1005
277 803
1 0 4 0 0 4096 0 3 0 0 9 3
529 954
808 954
808 747
7 4 4 0 0 8320 0 13 10 0 0 3
799 747
1005 747
1005 234
0 0 3 0 0 0 0 0 0 55 11 3
351 341
351 349
365 349
0 2 3 0 0 0 0 0 6 0 0 4
365 344
365 448
697 448
697 331
1 6 5 0 0 8320 0 9 8 0 0 5
970 236
970 297
491 297
491 320
468 320
2 0 6 0 0 8320 0 9 0 0 17 3
964 236
964 302
612 302
3 6 7 0 0 8320 0 9 6 0 0 3
958 236
958 322
752 322
3 1 8 0 0 4224 0 4 6 0 0 3
697 226
697 322
704 322
1 0 5 0 0 0 0 4 0 0 22 5
652 217
542 217
542 199
468 199
468 221
6 2 6 0 0 0 0 7 4 0 0 3
612 324
612 235
652 235
3 1 9 0 0 4224 0 5 7 0 0 3
531 229
531 324
564 324
2 5 10 0 0 8320 0 5 6 0 0 5
486 238
486 287
769 287
769 340
758 340
3 0 5 0 0 0 0 7 0 0 21 2
564 342
485 342
6 3 5 0 0 0 0 8 6 0 0 5
468 320
485 320
485 377
704 377
704 340
6 1 5 0 0 0 0 8 5 0 0 5
468 320
468 221
472 221
472 220
486 220
4 0 11 0 0 4096 0 8 0 0 25 4
444 368
444 383
448 383
448 391
4 0 11 0 0 4112 0 7 0 0 25 2
588 372
588 391
0 4 11 0 0 8320 0 0 6 26 0 4
409 344
409 391
728 391
728 370
0 3 11 0 0 0 0 0 8 27 0 5
409 326
409 344
409 344
409 338
420 338
1 1 11 0 0 0 0 1 8 0 0 6
333 267
409 267
409 326
409 326
409 320
420 320
2 0 3 0 0 0 0 7 0 0 11 3
557 333
554 333
554 448
1 0 2 0 0 8320 0 10 0 0 40 4
1023 234
1023 705
305 705
305 755
2 0 12 0 0 8320 0 10 0 0 38 4
1017 234
1017 710
472 710
472 757
3 7 13 0 0 4224 0 10 14 0 0 5
1011 234
1011 715
653 715
653 748
639 748
0 0 2 0 0 0 0 0 0 33 42 4
524 544
398 544
398 645
326 645
1 0 2 0 0 0 0 11 0 0 37 5
654 558
654 544
523 544
523 553
506 553
2 0 12 0 0 0 0 11 0 0 38 4
645 558
645 535
485 535
485 563
3 7 13 0 0 0 0 11 14 0 0 9
636 558
636 546
612 546
612 652
626 652
626 678
669 678
669 748
639 748
4 2 14 0 0 12416 0 11 13 0 0 6
645 603
645 655
718 655
718 743
751 743
751 747
0 1 2 0 0 0 0 0 17 42 0 5
326 624
430 624
430 553
507 553
507 563
2 7 12 0 0 0 0 17 15 0 0 4
489 563
477 563
477 757
468 757
1 6 15 0 0 8320 0 18 13 0 0 5
371 564
371 530
911 530
911 765
805 765
7 0 2 0 0 0 0 16 0 0 42 2
301 755
326 755
0 4 2 0 0 0 0 0 15 42 0 2
326 775
420 775
2 4 2 0 0 0 0 18 13 0 0 5
353 564
326 564
326 870
751 870
751 765
3 2 16 0 0 4224 0 17 14 0 0 3
498 608
498 748
591 748
3 2 17 0 0 4224 0 18 15 0 0 3
362 609
362 757
420 757
0 4 18 0 0 12288 0 0 16 46 0 4
227 755
234 755
234 773
253 773
0 2 18 0 0 4096 0 0 16 50 0 3
227 694
227 755
253 755
0 1 18 0 0 0 0 0 16 50 0 2
277 694
277 728
0 1 18 0 0 0 0 0 15 50 0 2
444 694
444 730
0 1 18 0 0 0 0 0 14 50 0 2
615 694
615 721
1 1 18 0 0 4224 0 2 13 0 0 3
191 694
775 694
775 720
3 0 19 0 0 8192 0 15 0 0 53 3
414 766
410 766
410 883
3 0 19 0 0 8192 0 14 0 0 53 3
585 757
577 757
577 883
0 3 19 0 0 8320 0 0 13 54 0 4
185 748
185 883
745 883
745 756
3 3 19 0 0 0 0 12 16 0 0 4
135 748
239 748
239 764
247 764
2
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 15
396 484 679 532
409 493 665 525
15 Circuito MOD-10
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
429 150 694 198
442 159 680 191
14 Circuito MOD-6
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
